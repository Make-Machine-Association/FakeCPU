module FakeCPU();

endmodule
